LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE VgaUtils IS
  CONSTANT COLOR_WHITE : STD_LOGIC_VECTOR := "111";
  CONSTANT COLOR_YELLOW : STD_LOGIC_VECTOR := "110";
  CONSTANT COLOR_PURPLE : STD_LOGIC_VECTOR := "101";
  CONSTANT COLOR_RED : STD_LOGIC_VECTOR := "100";
  CONSTANT COLOR_WATER : STD_LOGIC_VECTOR := "011";
  CONSTANT COLOR_GREEN : STD_LOGIC_VECTOR := "010";
  CONSTANT COLOR_BLUE : STD_LOGIC_VECTOR := "001";
  CONSTANT COLOR_BLACK : STD_LOGIC_VECTOR := "000";

  -- Timing values for 640x480@60Hz resolution
  -- http://tinyvga.com/vga-timing/640x480@60Hz
  CONSTANT H_SYNC_PULSE : INTEGER := 96;
  CONSTANT H_BACK_PORCH : INTEGER := 48;
  CONSTANT H_PIXELS : INTEGER := 640;
  CONSTANT H_FRONT_PORCH : INTEGER := 16;
  CONSTANT H_SYNC_POLARITY : STD_LOGIC := '0';

  CONSTANT V_SYNC_PULSE : INTEGER := 2;
  CONSTANT V_BACK_PORCH : INTEGER := 33;
  CONSTANT V_PIXELS : INTEGER := 480;
  CONSTANT V_FRONT_PORCH : INTEGER := 10;
  CONSTANT V_SYNC_POLARITY : STD_LOGIC := '0';

  -- Timing values for 800x600@72Hz resolution
  -- http://tinyvga.com/vga-timing/800x600@72Hz
  -- If using these timings, use the 50MHz clock directly instead of dividing by 2
  -- CONSTANT H_SYNC_PULSE : INTEGER := 120;
  -- CONSTANT H_BACK_PORCH : INTEGER := 64;
  -- CONSTANT H_PIXELS : INTEGER := 800;
  -- CONSTANT H_FRONT_PORCH : INTEGER := 56;
  -- CONSTANT H_SYNC_POLARITY : STD_LOGIC := '1';

  -- CONSTANT V_SYNC_PULSE : INTEGER := 6;
  -- CONSTANT V_BACK_PORCH : INTEGER := 23;
  -- CONSTANT V_PIXELS : INTEGER := 600;
  -- CONSTANT V_FRONT_PORCH : INTEGER := 37;
  -- CONSTANT V_SYNC_POLARITY : STD_LOGIC := '1';
END PACKAGE;

PACKAGE BODY VgaUtils IS
END VgaUtils;