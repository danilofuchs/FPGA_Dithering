LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY VgaOutput IS
    PORT (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC

    );
END ENTITY VgaOutput;

ARCHITECTURE rtl OF VgaOutput IS

BEGIN

END ARCHITECTURE;